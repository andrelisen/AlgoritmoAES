library verilog;
use verilog.vl_types.all;
entity memoria_chave_vlg_vec_tst is
end memoria_chave_vlg_vec_tst;
