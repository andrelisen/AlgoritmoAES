library verilog;
use verilog.vl_types.all;
entity AES_vlg_vec_tst is
end AES_vlg_vec_tst;
