library verilog;
use verilog.vl_types.all;
entity SubBytes_vlg_vec_tst is
end SubBytes_vlg_vec_tst;
