library verilog;
use verilog.vl_types.all;
entity memoria_sbox_vlg_vec_tst is
end memoria_sbox_vlg_vec_tst;
