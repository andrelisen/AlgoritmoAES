library verilog;
use verilog.vl_types.all;
entity ShiftRows is
    port(
        e0              : in     vl_logic_vector(7 downto 0);
        e1              : in     vl_logic_vector(7 downto 0);
        e2              : in     vl_logic_vector(7 downto 0);
        e3              : in     vl_logic_vector(7 downto 0);
        e4              : in     vl_logic_vector(7 downto 0);
        e5              : in     vl_logic_vector(7 downto 0);
        e6              : in     vl_logic_vector(7 downto 0);
        e7              : in     vl_logic_vector(7 downto 0);
        e8              : in     vl_logic_vector(7 downto 0);
        e9              : in     vl_logic_vector(7 downto 0);
        e10             : in     vl_logic_vector(7 downto 0);
        e11             : in     vl_logic_vector(7 downto 0);
        e12             : in     vl_logic_vector(7 downto 0);
        e13             : in     vl_logic_vector(7 downto 0);
        e14             : in     vl_logic_vector(7 downto 0);
        e15             : in     vl_logic_vector(7 downto 0);
        s0              : out    vl_logic_vector(7 downto 0);
        s1              : out    vl_logic_vector(7 downto 0);
        s2              : out    vl_logic_vector(7 downto 0);
        s3              : out    vl_logic_vector(7 downto 0);
        s4              : out    vl_logic_vector(7 downto 0);
        s5              : out    vl_logic_vector(7 downto 0);
        s6              : out    vl_logic_vector(7 downto 0);
        s7              : out    vl_logic_vector(7 downto 0);
        s8              : out    vl_logic_vector(7 downto 0);
        s9              : out    vl_logic_vector(7 downto 0);
        s10             : out    vl_logic_vector(7 downto 0);
        s11             : out    vl_logic_vector(7 downto 0);
        s12             : out    vl_logic_vector(7 downto 0);
        s13             : out    vl_logic_vector(7 downto 0);
        s14             : out    vl_logic_vector(7 downto 0);
        s15             : out    vl_logic_vector(7 downto 0)
    );
end ShiftRows;
