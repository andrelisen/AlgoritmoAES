
library ieee;
use ieee.std_logic_1164.all;

entity controle_AES is
    port (
			--SINAL DE ENTRADA PARA A MAQ DE ESTADOS FUNCIONAR
			clock : in std_logic;
			reset : in std_logic;
			--SINAIS DE SAÃDA CALCULADOS PELA MAQ DE ESTADOS
			--Sinal de enable
			Enable_registradoresA	:	out std_logic;	--Inicializa 8 registradores
			Enable_registradoresB	:	out std_logic;	--Inicializa 8 registradores
			Enable_registradoresC	:	out std_logic;	--Inicializa 8 registradores
			Enable_registradoresD	:	out std_logic;	--Inicializa 8 registradores
			Enable_Add 					:	out std_logic;
			Enable_SubBytes			:  out std_logic;
			Enable_ShiftRows			:  out std_logic;
			Enable_Mix					:  out std_logic;
			Enable_SubChave			:  out std_logic;
		--Seletores
			Sel_EntradaAddTxt 		: out std_logic_vector(1 downto 0); -- entrada mux add txt
			Sel_EntradaAddKey 		: out std_logic;						  -- entrada mux add sub chave
			Sel_EntradaSubChave 		: out std_logic;
			Sel_rcon						: out std_logic_vector(3 downto 0)
    );
end entity;

architecture implementa of controle_AES is

   type type_state is 
		(state1, state2, state3, state4, state5, state6, state7, state8, state9, 
			state10, state11, state12, state13, state14, state15, state16, state17, state18, state19, state20,
			state21, state22, state23, state24, state25, state26, state27, state28, state29, state30,
			state31, state32, state33, state34, state35,state36, state37, state38, state39, state40, state41, state42,
			state43, state44, state45, state46, state47, state48, state49,state50 ,state51, state52, state53, state54
	);

	signal state: type_state;

begin

	 process (clock,reset)
    begin
        if (reset='1') then -- vai para o estado inicial sem borda de clock
            state <= state1;
        elsif(rising_edge(clock)) then
            case state is
					 when state1 =>
						  state <= state2;
					 when state2 =>
						  state <= state3;
					 when state3 =>
						  state <= state4;
					 when state4 =>
							state <= state5;
					 when state5 =>
							state <= state6;
					 when state6 =>
							state <= state7;
					 when state7 =>
						  state <= state8;
					 when state8 =>
						  state <= state9;
					 when state9 =>
						  state <= state10;
					 when state10 =>
						  state <= state11;
					 when state11 =>
						  state <= state12;
					 when state12 =>
						  state <= state13;
					 when state13 =>
						  state <= state14;
					 when state14 =>
						  state <= state15;
					 when state15 =>
						  state <= state16;
					 when state16 =>
							state <= state17;
					 when state17 =>
							state <= state18;
					 when state18 =>
							state <= state19;
					 when state19 =>
							state <= state20;
					 when state20 =>
						  state <= state21;
					 when state21 =>
							state <= state22;
					 when state22 =>
							state <= state23;
					 when state23 =>
							state <= state24;
					 when state24 =>
							state <= state25;
					 when state25 => 
							state <= state26;
					 when state26 => 
							state <= state27;
					 when state27 => 
							state <= state28;
					when state28 => 
							state <= state29;
					when state29 => 
							state <= state30;
					when state30 => 
							state <= state31;
					when state31 => 
							state <= state32;
					when state32 => 
							state <= state33;
					when state33 => 
							state <= state34;
					when state34 => 
							state <= state35;
					when state35 => 
							state <= state36;
					when state36 => 
							state <= state37;
					when state37 => 
							state <= state38;
					when state38 => 
							state <= state39;
					when state39 => 
							state <= state40;
					when state40 => 
							state <= state41;
					when state41 => 
							state <= state42;
					when state42 => 
							state <= state43;
					when state43 => 
							state <= state44;
					when state44 => 
							state <= state45;
					when state45 => 
							state <= state46;
					when state46 => 
							state <= state47;
					when state47 => 
							state <= state48;
					when state48 => 
							state <= state49;
					when state49 => 
							state <= state50;
					when state50 => 
							state <= state51;
					when state51 => 
							state <= state52;
					when state52 => 
							state <= state53;
					when state53 => 
							state <= state54;
					 when others => 
							state <= state54;
            end case;
        end if;
    end process;

    process (state) --bloco combinacional: saÃ­das sÃ£o calculadas em funÃ§Ã£o do estado atual do controle.
    begin			  
		case state is
			 when state1 => -- INICIALIZA REG
				Enable_registradoresA	<= '1';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
			 when state2 => -- INICIALIZA REG
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '1';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
			 when state3 => -- INICIALIZA REG
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '1';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
			 when state4 => -- INICIALIZA REG
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '1';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
			 when state5 => -- ADD KEY COM CHAVE INICIAL 1
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
			 when state6 => --calculo sub chave1
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "00";
				Sel_EntradaAddKey 		<= '1';
				Sel_EntradaSubChave 		<='1';
				Sel_rcon						<="0001";
				when state7 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0010";
				when state8 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0010";
				when state9 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0010";
				when state10 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0010";
				when state11 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0010";
				when state12 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0011";
				when state13 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0011";
				when state14 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0011";
				when state15 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0011";
				when state16 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0011";
				when state17 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0100";
				when state18 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0100";
				when state19 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0100";
				when state20 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0100";
				when state21 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0100";
				when state22 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0101";
				when state23 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0101";
				when state24 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0101";
				when state25 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0101";
				when state26 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0101";
				when state27 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0110";
				when state28 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0110";
				when state29 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0110";
				when state30 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0110";
				when state31 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0110";
				when state32 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0111";
				when state33 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0111";
				when state34 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0111";
				when state35 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0111";
				when state36 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="0111";
				when state37 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1000";
				when state38 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1000";
				when state39 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1000";
				when state40 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1000";
				when state41 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1000";
				when state42 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1001";
				when state43 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1001";
				when state44 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1001";
				when state45 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1001";
				when state46 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1001";
				
				when state47 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state48 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state49 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '1';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state50 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state51 => --calculo sub chave
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '1';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				
				when state52 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '1';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state53 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '0';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '1';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "01";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				when state54 => 
				Enable_registradoresA	<= '0';
				Enable_registradoresB	<= '0';
				Enable_registradoresC	<= '0';
				Enable_registradoresD	<= '0';
				Enable_Add 					<= '1';
				Enable_SubBytes			<= '0';
				Enable_ShiftRows			<= '0';
				Enable_Mix					<= '0';
				Enable_SubChave			<= '0';
				Sel_EntradaAddTxt 		<= "10";
				Sel_EntradaAddKey 		<= '0';
				Sel_EntradaSubChave 		<='0';
				Sel_rcon						<="1010";
				
 		end case;
    end process;          
	 
end implementa;
