library verilog;
use verilog.vl_types.all;
entity SubChave_vlg_vec_tst is
end SubChave_vlg_vec_tst;
