library verilog;
use verilog.vl_types.all;
entity ShiftRows_vlg_vec_tst is
end ShiftRows_vlg_vec_tst;
