library verilog;
use verilog.vl_types.all;
entity MixColumns_vlg_vec_tst is
end MixColumns_vlg_vec_tst;
