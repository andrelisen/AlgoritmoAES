library verilog;
use verilog.vl_types.all;
entity Conecta_topo_vlg_vec_tst is
end Conecta_topo_vlg_vec_tst;
