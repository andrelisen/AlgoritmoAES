library verilog;
use verilog.vl_types.all;
entity AES_topo_vlg_vec_tst is
end AES_topo_vlg_vec_tst;
