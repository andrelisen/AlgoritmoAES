library verilog;
use verilog.vl_types.all;
entity SubChave_vlg_check_tst is
    port(
        n0              : in     vl_logic_vector(7 downto 0);
        n1              : in     vl_logic_vector(7 downto 0);
        n2              : in     vl_logic_vector(7 downto 0);
        n3              : in     vl_logic_vector(7 downto 0);
        n4              : in     vl_logic_vector(7 downto 0);
        n5              : in     vl_logic_vector(7 downto 0);
        n6              : in     vl_logic_vector(7 downto 0);
        n7              : in     vl_logic_vector(7 downto 0);
        n8              : in     vl_logic_vector(7 downto 0);
        n9              : in     vl_logic_vector(7 downto 0);
        n10             : in     vl_logic_vector(7 downto 0);
        n11             : in     vl_logic_vector(7 downto 0);
        n12             : in     vl_logic_vector(7 downto 0);
        n13             : in     vl_logic_vector(7 downto 0);
        n14             : in     vl_logic_vector(7 downto 0);
        n15             : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end SubChave_vlg_check_tst;
