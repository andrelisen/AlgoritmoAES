library verilog;
use verilog.vl_types.all;
entity Conecta_topo_vlg_check_tst is
    port(
        out0Add_top     : in     vl_logic_vector(7 downto 0);
        out1Add_top     : in     vl_logic_vector(7 downto 0);
        out2Add_top     : in     vl_logic_vector(7 downto 0);
        out3Add_top     : in     vl_logic_vector(7 downto 0);
        out4Add_top     : in     vl_logic_vector(7 downto 0);
        out5Add_top     : in     vl_logic_vector(7 downto 0);
        out6Add_top     : in     vl_logic_vector(7 downto 0);
        out7Add_top     : in     vl_logic_vector(7 downto 0);
        out8Add_top     : in     vl_logic_vector(7 downto 0);
        out9Add_top     : in     vl_logic_vector(7 downto 0);
        out10Add_top    : in     vl_logic_vector(7 downto 0);
        out11Add_top    : in     vl_logic_vector(7 downto 0);
        out12Add_top    : in     vl_logic_vector(7 downto 0);
        out13Add_top    : in     vl_logic_vector(7 downto 0);
        out14Add_top    : in     vl_logic_vector(7 downto 0);
        out15Add_top    : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Conecta_topo_vlg_check_tst;
