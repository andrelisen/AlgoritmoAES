library verilog;
use verilog.vl_types.all;
entity Mux10p1_vlg_vec_tst is
end Mux10p1_vlg_vec_tst;
